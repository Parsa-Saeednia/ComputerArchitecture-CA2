module Alu();
    
    
endmodule