`timescale 1ns/1ns
module Extend(imm, immSrc, immExt);
    input [31:7] imm;
    input [1:0] immSrc;
    output [31:0] immExt;
    
    
endmodule