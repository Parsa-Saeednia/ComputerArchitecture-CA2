module Datapath();
    
    
endmodule